module top_module(
    output zero
);// Module body starts after semicolon
//Left this blank since not assigning a value will lead to 0, in simulation
  assign zero = 1'b0;
endmodule
