module top_module( output one );

// Insert your code here
    assign one = 1;
    //my solution is 1, suggested is 1'b1

endmodule
